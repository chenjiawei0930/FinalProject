module dodge(output reg [7:0] DATA_R, DATA_G, DATA_B,output reg [2:0] COMM,output reg EN, input CLK, clear, Left, Right, Up,Down,
                                                                                    output reg [3:0] Life,
									output reg [6:0] d7_1,    
								                    output reg [1:0] COMM_CLK)	;															  

reg [7:0] plate [7:0];
reg [7:0] people [7:0];
reg [6:0] seg1, seg2;
reg [3:0] bcd_s,bcd_m;
segment7 S0(bcd_s, A0,B0,C0,D0,E0,F0,G0);
segment7 S1(bcd_m, A1,B1,C1,D1,E1,F1,G1);
divfreq div0(CLK, CLK_div);
divfreq1(CLK, CLK_time);
divfreq2 div2(CLK, CLK_mv);
reg [2:0] random01, random02, random03,random04,random05, r, r1, r2,r3,r4;
reg left, right,up,down;
integer a,b,c,d,e,count,line,row,touch,count1;
initial
begin 
a=0;
b=0;
c=0;
d=0;
e=7;
line = 3;
row=6;
touch=0;
bcd_m = 0;
bcd_s = 0;
random01 = (5*random01 + 3)%16;
			r = random01 % 8;
random02 = (5*(random02+1) + 3)%16;
        r1 = random02 % 8;
random03= (5*(random03+2) + 3)%16;
			r2 = random03 % 8;
random04= (5*(random04+3) + 3)%16;
			r3 = random04 % 8;
random05= (5*(random05+4) + 3)%16;
			r4 = random05 % 8;			
			DATA_R = 8'b11111111;
			DATA_G = 8'b11111111;
			DATA_B = 8'b11111111;
			plate[0] = 8'b11111111;
			plate[1] = 8'b11111111;
			plate[2] = 8'b11111111;
			plate[3] = 8'b11111111;
			plate[4] = 8'b11111111;
			plate[5] = 8'b11111111;
			plate[6] = 8'b11111111;
			plate[7] = 8'b11111111;
			people[0] = 8'b11111111;
			people[1] = 8'b11111111;
			people[2] = 8'b11111111;
			people[3] = 8'b00111111;
			people[4] = 8'b11111111;
			people[5] = 8'b11111111;
			people[6] = 8'b11111111;
			people[7] = 8'b11111111;
			count1=0;
		
end 

always@(posedge CLK_div)
	begin
		seg1[0] = A0;
		seg1[1] = B0;
		seg1[2] = C0;
		seg1[3] = D0;
		seg1[4] = E0;
		seg1[5] = F0;
		seg1[6] = G0;
		
		seg2[0] = A1;
		seg2[1] = B1;
		seg2[2] = C1;
		seg2[3] = D1;
		seg2[4] = E1;
		seg2[5] = F1;
		seg2[6] = G1;
		
		if(count1 == 0)
			begin
				d7_1 <= seg1;
				COMM_CLK[1] <= 1'b1;
				COMM_CLK[0] <= 1'b0;
				count1 <= 1'b1;
			end
		else if(count1 == 1)
			begin
				d7_1 <= seg2;
				COMM_CLK[1] <= 1'b0;
				COMM_CLK[0] <= 1'b1;
				count1 <= 1'b0;
			end
		
		


	end
always@(posedge CLK_time, posedge clear)
	begin
		if(clear)
			begin
				bcd_m = 3'b0;
				bcd_s = 4'b0;
			end
		else
			begin
				if(touch < 3)
					begin
						if(bcd_s >= 9)
							begin
								bcd_s <= 0;
								bcd_m <= bcd_m + 1;
							end
						else
							bcd_s <= bcd_s + 1;
						if(bcd_m >= 9) bcd_m <= 0;
					end
			end
	end


	always@(posedge CLK_div)
	begin
		if(count >= 7)
			count <= 0;
		else
		count <= count + 1;
		
		COMM =count;
		EN = 1'b1;
		if(touch < 4)
			begin
				DATA_G <= plate[count];
				DATA_R <= people[count];
				if(touch == 0)
					Life <= 4'b1111;
				else if(touch == 1)
					Life <= 4'b1110;
				else if(touch == 2)
					Life <= 4'b1100;
				else if(touch == 3)
					Life <= 4'b1000;	
			end
		else
			begin
				DATA_R <= plate[count];
				DATA_G <= 8'b11111111;
				Life <= 4'b0000;
			end
			
	
		
				
		
	end
//遊戲
always@(posedge CLK_mv)
	begin
	    right = Right;
		 left=Left;
		 up=Up;
		 down=Down;
		if(clear==1)
	     begin
		         touch = 0;
					line = 3;
					a = 0;
					b = 0;
					c = 0;
					d=3;
					e=7;
					row=6;
					random01 = (5*random01 + 3)%16;
					r = random01 % 8;
					random02 = (5*(random02+1) + 3)%16;
					r1 = random02 % 8;
					random03= (5*(random03+2) + 3)%16;
					r2 = random03 % 8;
					random04= (5*(random04+2) + 3)%16;
			     r3 = random04 % 8;
             random05= (5*(random05+2) + 3)%16;
			      r4 = random05 % 8;			
					plate[0] = 8'b11111111;
					plate[1] = 8'b11111111;
					plate[2] = 8'b11111111;
					plate[3] = 8'b11111111;
					plate[4] = 8'b11111111;
					plate[5] = 8'b11111111;
					plate[6] = 8'b11111111;
					plate[7] = 8'b11111111;
					people[0] = 8'b11111111;
					people[1] = 8'b11111111;
					people[2] = 8'b11111111;
					people[3] = 8'b00111111;
					people[4] = 8'b11111111;
					people[5] = 8'b11111111;
					people[6] = 8'b11111111;
					people[7] = 8'b11111111;
			end
  if(touch < 4)
	begin	
	//fall object 1
		/*if(a == 0)
					begin
						plate[r][a] = 1'b0;
						a = a+1;
					end
				else if (a > 0 && a <= 7)
						begin
							plate[r][a-1] = 1'b1;
							plate[r][a] = 1'b0;
							a = a+1;
						end
				else if(a == 8) 
					begin
						plate[r][a-1] = 1'b1;
						random01 = (5*random01 + 3)%16;
						r = random01 % 8;
						a = 0;
		          end
		*/
			//fall object 2
			if(b == 0)
					begin
						plate[r1][b] = 1'b0;
						b = b+1;
					end
				else if (b > 0 && b <= 7)
					begin
						plate[r1][b-1] = 1'b1;
						plate[r1][b] = 1'b0;
						b = b+1;
					end
				else if(b == 8) 
					begin
						plate[r1][b-1] = 1'b1;
						random02 = (5*(random02+1) + 3)%16;
						r1 = random02 % 8;
						b = 0;
					end	
					
			if(c == 0)
					begin
						plate[r2][c] = 1'b0;
						c = c+1;
					end
				else if (c > 0 && c <= 7)
					begin
						plate[r2][c-1] = 1'b1;
						plate[r2][c] = 1'b0;
						c = c+1;
					end
				else if(c == 8) 
					begin
						plate[r2][c-1] = 1'b1;
						random03= (5*(random03+2) + 3)%16;
						r2 = random03 % 8;
						c = 0;
					end
				
		if (d==0)
              begin
				plate[d][r3]=1'b0;
		       d=d+1;
			    end
			else if (d>0 && d<=7)
	        begin 
			       plate[d-1][r3]=1'b1;
				    plate[d][r3]=1'b0;
				    d=d+1;	 
				end	
			else if(d == 8) 
					begin
						plate[d-1][r3] = 1'b1;
						random04= (5*(random04+2) + 3)%16;
						r3=random04 % 8;
						d =0;
					end	
					
		if (e==7)
             begin
				plate[e][r4]=1'b0;
		       e=e-1;
			    end
			else if (e>0 && e<7)
	        begin 
			       plate[e+1][r4]=1'b1;
				    plate[e][r4]=1'b0;
				    e=e-1;	 
				end	
			else if(e == -1) 
					begin
						plate[e+1][r4] = 1'b1;
						random05= (5*(random05+4) + 3)%16;
						r4=random05 % 8;
						e =7;
			end				
		//pepole move
 if(right == 1 || left ==1 )
	begin
		if((right == 1) && (line != 7))
					begin
						people[line][row] = 1'b1;
						people[line][row+1] = 1'b1;
						line = line + 1;
					end
		if((left == 1) && (line != 0))
					begin
						people[line][row] = 1'b1;
						people[line][row+1] = 1'b1;
						line = line - 1;
					end
		 people[line][row] = 1'b0;
		 people[line][row+1] = 1'b0;
	end	 
else if (up == 1 || down == 1)
  begin 
		if( (up == 1) && (row != 0)) 
           begin	
			   people[line][row+1] = 1'b1;
			   row =row -1;
				people[line][row] = 1'b0;	
			  end	
		if(  (down == 1) && row!= 6 )	  
       begin	
			   people[line][row] = 1'b1;
			  row =row +1;
				people[line][row+1] = 1'b0;	
		 end
 	
	end	
	   
			  
		 if(plate[line][row] == 0)
					begin
						touch = touch + 1;
						plate[r][row] = 1'b1;
						
						plate[r1][row] = 1'b1;
						
						plate[r2][row] = 1'b1;
						
						plate[r3][row] = 1'b1;
						plate[r4][row] = 1'b1;
						
						a = 8;
						b = 8;
						c = 8;
						d = 8;
						e = -1;
					end
		else if (plate[line][row+1] == 0)
			begin
						touch = touch + 1;
												
						plate[r][row+1] = 1'b1;
						
						plate[r1][row+1] = 1'b1;
						
						plate[r2][row+1] = 1'b1;
						plate[r3][row+1] = 1'b1;
						
						plate[r4][row+1] = 1'b1;
						a = 8;
						b = 8;
						c = 8;
						d = 8;
						e = -1;
						
				end
	end	
		else
			begin
				plate[0] = 8'b01101110;
				plate[1] = 8'b10110101;                      
            plate[2] = 8'b10111011;
				plate[3] = 8'b10111111;
				plate[4] = 8'b10111111;
				plate[5] = 8'b10111011;
				plate[6] = 8'b10110101;
				plate[7] = 8'b01101110;
			end			
		
						
					
end
endmodule





module segment7(input [0:3] a, output A,B,C,D,E,F,G);


	
	assign A = ~(a[0]&~a[1]&~a[2] | ~a[0]&a[2] | ~a[1]&~a[2]&~a[3] | ~a[0]&a[1]&a[3]),
	       B = ~(~a[0]&~a[1] | ~a[1]&~a[2] | ~a[0]&~a[2]&~a[3] | ~a[0]&a[2]&a[3]),
			 C = ~(~a[0]&a[1] | ~a[1]&~a[2] | ~a[0]&a[3]),
			 D = ~(a[0]&~a[1]&~a[2] | ~a[0]&~a[1]&a[2] | ~a[0]&a[2]&~a[3] | ~a[0]&a[1]&~a[2]&a[3] | ~a[1]&~a[2]&~a[3]),
			 E = ~(~a[1]&~a[2]&~a[3] | ~a[0]&a[2]&~a[3]),
			 F = ~(~a[0]&a[1]&~a[2] | ~a[0]&a[1]&~a[3] | a[0]&~a[1]&~a[2] | ~a[1]&~a[2]&~a[3]),
			 G = ~(a[0]&~a[1]&~a[2] | ~a[0]&~a[1]&a[2] | ~a[0]&a[1]&~a[2] | ~a[0]&a[2]&~a[3]);
			 
endmodule





//計時除頻器
module divfreq1(input CLK, output reg CLK_time);
  reg [25:0] Count;
  initial
    begin
      CLK_time = 0;
	 end	
		
  always @(posedge CLK)
    begin
      if(Count > 25000000)
        begin
          Count <= 25'b0;
          CLK_time <= ~CLK_time;
        end
      else
        Count <= Count + 1'b1;
    end
endmodule 











//視覺暫留除頻器
module divfreq(input CLK, output reg CLK_div);
  reg [24:0] Count;
  always @(posedge CLK)
    begin
      if(Count > 10000)
        begin
          Count <= 25'b0;
          CLK_div <= ~CLK_div;
        end
      else
        Count <= Count + 1'b1;
    end
endmodule

//掉落物&人物移動除頻器
module divfreq2(input CLK, output reg CLK_mv);
  reg [35:0] Count;
  initial
    begin
      CLK_mv = 0;
	 end	
		
  always @(posedge CLK)
    begin
      if(Count > 3500000)
        begin
          Count <= 35'b0;
          CLK_mv <= ~CLK_mv;
        end
      else
        Count <= Count + 1'b1;
    end
endmodule 
